`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/26/2022 11:17:12 PM
// Design Name: 
// Module Name: fpga_wrap
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fpga_wrap(
    input logic CLK100, 
    input logic [15:0] SW, 
    output logic [15:0] LED, 
    output logic [7:0] AN,

    );
endmodule
